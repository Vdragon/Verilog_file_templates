//include guard
`ifndef 
	`define 
	// 時間相關設定
	`timescale 1ns / 100ps

	/* 模組名稱 | Module Name
				
		 著作權宣告 | Copyright Declaration
				copyright 2012 林博仁(pika1021@gmail.com) */
	module ();
	//port 輸出輸入宣告
	output ;
	input ;

	//port 類型宣告
	reg ;
	wire ;

	endmodule
`endif