/* 模組名稱：
   著作權宣告：copyright 2012 林博仁(pika1021@gmail.com)
   */
`timescale 1ns / 100ps

module ();
  output
  input
endmodule
